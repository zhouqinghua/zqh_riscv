#defaultvalue x|z|0|1|random|random seed_value
#instance instance_hierarchical_name [x|z|0|1|random|
#random seed_value]
#tree instance_hierarchical_name depth [x|z|0|1|random|
#random seed_value]
#module module_name [x|z|0|1|random|random seed_value]
#modtree module_name depth [x|z|0|1|random|
#random seed_value]

defaultvalue random
tree top.test_harness.dut 0 random
